module testModule (
    input d,
    output o
);
    assign o = !d;

endmodule


